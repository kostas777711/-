** Profile: "SCHEMATIC1-lag filter"  [ D:\ORCAD\WORKS DIPLOMATIKHS\lag filter-SCHEMATIC1-lag filter.sim ] 

** Creating circuit file "lag filter-SCHEMATIC1-lag filter.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\ORCAD\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 20ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\lag filter-SCHEMATIC1.net" 


.END
